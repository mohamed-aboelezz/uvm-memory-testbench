`include "uvm_macros.svh"
package tb_pkg;
import uvm_pkg::*;

`include "package/my_sequence_item.sv"
`include "package/my_sequence.sv"
`include "package/my_driver.sv"
`include "package/my_sequencer.sv"
`include "package/my_monitor.sv"
`include "package/my_subscriber.sv"
`include "package/my_scoreboard.sv"
`include "package/my_agent.sv"
`include "package/my_env.sv"
`include "package/my_test.sv"

endpackage